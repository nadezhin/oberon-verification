`timescale 1ns / 1ps
module BUFG(input I, output O);
assign O = I;
endmodule
