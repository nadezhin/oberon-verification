`timescale 1ns / 1ps
module IBUFG(input I, output O);
assign O = I;
endmodule
